.TITLE Hugo Frisk Op-Amp


.SUBCKT opAmp vdd vddOutputStage vss vssOutputStage inputP inputN output
.INCLUDE irlml2246trpbf.spi	$ P-channel signal MOSFET - drain, gate, source
.INCLUDE irlml6346trpbf.spi	$ N-channel signal MOSFET - drain, gate, source
.INCLUDE irf5305.spi		$ P-channel power MOSFET - drain, gate, source
.INCLUDE irfz48vs.spi 		$ N-channel power MOSFET - drain, gate, source

* Current mirror for tail current and biasing in intermediate stage
R11 vdd ISet 10k
X11 ISet ISet vss irlml6346trpbf

* Input pair
X21 inDrainP inputP tail irlml6346trpbf
X22 inDrainN inputN tail irlml6346trpbf 

* Tail
X23 tail ISet vss irlml6346trpbf

* Current mirror for input pair
X24 inDrainP inDrainP vdd irlml2246trpbf
X25 inDrainN inDrainP vdd irlml2246trpbf

* Intermediate stage
X31 outputPChGate inDrainN vdd irlml2246trpbf
C31 inDrainN outputPChGate 90p $ Compensation capacitor
R32 outputPChGate outputNChGate 5k
X32 outputNChGate ISet vss irlml6346trpbf

* Output stage
X41 output outputPChGate vddOutputStage irf5305
X42 output outputNChGate vssOutputStage IRFZ48VS 

.ENDS

X1 vdd vddOutputStage vss vssOutputStage in feedback out opAmp

* Power supply
VP vdd 0 DC 5	$ Positive rail
VN 0 vss DC 5	$ Negative rail
VPOutputStage vddOutputStage 0 DC 5 $ Seperate positive rail for output stage in order the mesure its current
VNOutputStage 0 vssOutputStage DC 5 $ Seperate negative rail for output stage in order the mesure its current

* Test setup
VIn in 0 DC 0 AC 10u SIN(0 100m 100 0 0 90) $ PULSE(-5 5 0 20m 20m 1 1) -550u offset for 0v intermediate
R1 out feedback 9k
R2 feedback 0 1k


.CONTROL
TRAN 100u 20m
PLOT in out XLIMIT 0 20m YLIMIT -5 5
PLOT out/in VS in XLIMIT -30m 30m

SET UNITS = degrees
AC DEC 10 1 1MEG
LET gain = V(out)/V(in)
PLOT DB(gain) XLIMIT 1 1MEG
PLOT CPH(out) XLIMIT 1 1MEG YLIMIT -360 0 YDELTA 45
MEAS AC maxGain MAX VDB(gain) FROM=1 TO=1MEG
.ENDC

.END
