.TITLE Hugo Frisk Op-Amp


.SUBCKT opAmp vdd vss inputP inputN output
.INCLUDE irlml2246trpbf.spi	$ P-channel signal MOSFET - drain, gate, source
.INCLUDE irlml6346trpbf.spi	$ N-channel signal MOSFET - drain, gate, source
.INCLUDE irf5305.spi		$ P-channel power MOSFET - drain, gate, source
.INCLUDE irfz48vs.spi 		$ N-channel power MOSFET - drain, gate, source

* Current mirror for tail current and biasing in intermediate stage
R11 vdd ISet 10k
X11 ISet ISet vss irlml6346trpbf

* Input pair
X21 inDrainP inputP tail irlml6346trpbf
X22 inDrainN inputN tail irlml6346trpbf 

* Tail
X23 tail ISet vss irlml6346trpbf

* Current mirror for input pair
X24 inDrainP inDrainP vdd irlml2246trpbf
X25 inDrainN inDrainP vdd irlml2246trpbf

* Intermediate stage
X31 outputPChGate inDrainN vdd irlml2246trpbf
R31 outputPChGate outputNChGate 4k
X32 outputNChGate ISet vss irlml6346trpbf

* Output stage
X41 output outputPChGate vdd irf5305
X42 output outputNChGate vss IRFZ48VS 

.ENDS

X1 vdd vss in 0 out opAmp

* Power supply
VP vdd 0 DC 5	$ Positive rail
VN 0 vss 5	$ Negative rail

* Test setup
VDiff in 0 SIN(0 100n 100 0 0 0)
* R1 out 0 100

.CONTROL
TRAN 100u 20m
PLOT in XLIMIT 0 20m
PLOT out XLIMIT 0 20m
PLOT X1.inDrainN XLIMIT 0 20m
PLOT X1.outputPChGate X1.outputNChGate XLIMIT 0 20m
.ENDC

.END
